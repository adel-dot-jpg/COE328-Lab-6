library verilog;
use verilog.vl_types.all;
entity lab6_Part3_vlg_vec_tst is
end lab6_Part3_vlg_vec_tst;
