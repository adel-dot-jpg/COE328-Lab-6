library ieee;
use ieee.std_logic_1164.all;

entity reg1 is
	port (
		A : in std_logic_vector(7 downto 0);
		res, clk : in std_logic;
		Q : out std_logic_vector(7 downto 0)
	);
end reg1;

architecture behavior of reg1 is
begin
	process(res, clk)
	begin
		if res = '1' then
			Q <= "00000000";
		elsif (clk'event and clk = '1') then
			Q <= A;
		end if;
	end process;
end behavior;