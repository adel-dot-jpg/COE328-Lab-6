LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_signed.all;

ENTITY signed_seg7 IS
PORT (
  bcd      : IN  STD_LOGIC_VECTOR(3 DOWNTO 0); -- signed input
  leds_mag : OUT STD_LOGIC_VECTOR(1 TO 7);     -- magnitude display
  leds_sign: OUT STD_LOGIC_VECTOR(1 TO 7)      -- sign display
);
END signed_seg7;

ARCHITECTURE Behavior OF signed_seg7 IS
  SIGNAL magnitude : STD_LOGIC_VECTOR(3 DOWNTO 0);
BEGIN
  PROCESS (bcd)
  BEGIN
    -- Sign logic
    IF bcd(3) = '1' THEN  -- Negative number
      leds_sign <= "0000001";  -- Dash (only g is ON)
      magnitude <= NOT(bcd) + 1;  -- Two's complement to get magnitude
    ELSE
      leds_sign <= "0000000";  -- No segments ON
      magnitude <= bcd;
    END IF;

    -- Magnitude to 7-seg
    CASE magnitude IS
      WHEN "0000" => leds_mag <= "1111110";  -- 0
      WHEN "0001" => leds_mag <= "0110000";  -- 1
      WHEN "0010" => leds_mag <= "1101101";  -- 2
      WHEN "0011" => leds_mag <= "1111001";  -- 3
      WHEN "0100" => leds_mag <= "0110011";  -- 4
      WHEN "0101" => leds_mag <= "1011011";  -- 5
      WHEN "0110" => leds_mag <= "1011111";  -- 6
      WHEN "0111" => leds_mag <= "1110000";  -- 7
      WHEN "1000" => leds_mag <= "1111111";  -- 8
      WHEN "1001" => leds_mag <= "1111011";  -- 9
      WHEN OTHERS => leds_mag <= "0000000";  -- off state? error state??
    END CASE;
  END PROCESS;
END Behavior;
